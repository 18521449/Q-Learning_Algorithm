module Register 
	#(	parameter WIDTH = 128)
	(	input valid_in,
		input clk,
		input [WIDTH-1:0] in,
		output [WIDTH-1:0] out, 
		output reg valid_out
	);

endmodule
